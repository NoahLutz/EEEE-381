** Profile: "SCHEMATIC1-differential_gain"  [ E:\Electronics 1 Lab\lab4\prelab\lab4_prelab-PSpiceFiles\SCHEMATIC1\differential_gain.sim ] 

** Creating circuit file "differential_gain.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.INC "../../../spice.txt" 
* From [PSPICE NETLIST] section of C:\Users\cnl9674\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
